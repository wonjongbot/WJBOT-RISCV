package wjbot_riscv;
	string proj_root = "/home/wonjongbot/WJBOT-RISCV/";
endpackage